netcdf tt {
dimensions:
	nele = xxxx ;
	node = xxxx ;
	siglay = 30 ;
	siglev = 31 ;
	three = 3 ;
	time = UNLIMITED ; // (1 currently)
	DateStrLen = 26 ;
variables:
	float x(node) ;
		x:long_name = "nodal x-coordinate" ;
		x:units = "meters" ;
	float y(node) ;
		y:long_name = "nodal y-coordinate" ;
		y:units = "meters" ;
	float lon(node) ;
		lon:long_name = "nodal longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	float lat(node) ;
		lat:long_name = "nodal latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	float xc(nele) ;
		xc:long_name = "zonal x-coordinate" ;
		xc:units = "meters" ;
	float yc(nele) ;
		yc:long_name = "zonal y-coordinate" ;
		yc:units = "meters" ;
	float lonc(nele) ;
		lonc:long_name = "zonal longitude" ;
		lonc:standard_name = "longitude" ;
		lonc:units = "degrees_east" ;
	float latc(nele) ;
		latc:long_name = "zonal latitude" ;
		latc:standard_name = "latitude" ;
		latc:units = "degrees_north" ;
	float siglay(siglay, node) ;
		siglay:long_name = "Sigma Layers" ;
		siglay:standard_name = "ocean_sigma/general_coordinate" ;
		siglay:positive = "up" ;
		siglay:valid_min = -1.f ;
		siglay:valid_max = 0.f ;
		siglay:formula_terms = "sigma: siglay eta: zeta depth: h" ;
	float siglev(siglev, node) ;
		siglev:long_name = "Sigma Levels" ;
		siglev:standard_name = "ocean_sigma/general_coordinate" ;
		siglev:positive = "up" ;
		siglev:valid_min = -1.f ;
		siglev:valid_max = 0.f ;
		siglev:formula_terms = "sigma:siglay eta: zeta depth: h" ;
	float h(node) ;
		h:long_name = "Bathymetry" ;
		h:standard_name = "sea_floor_depth_below_geoid" ;
		h:units = "m" ;
		h:positive = "down" ;
		h:grid = "Bathymetry_Mesh" ;
		h:coordinates = "x y" ;
		h:type = "data" ;
	int nv(three, nele) ;
		nv:long_name = "nodes surrounding element" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 1858-11-17 00:00:00" ;
		time:format = "modified julian day (MJD)" ;
		time:time_zone = "UTC" ;
	char Times(time, DateStrLen) ;
		Times:time_zone = "UTC" ;
	float zeta(time, node) ;
		zeta:long_name = "Water Surface Elevation" ;
		zeta:units = "meters" ;
		zeta:positive = "up" ;
		zeta:standard_name = "sea_surface_height_above_geoid" ;
		zeta:grid = "TWOD_Mesh" ;
		zeta:coordinates = "x y" ;
		zeta:type = "data" ;
	float u(time, siglay, nele) ;
		u:long_name = "Eastward Water Velocity" ;
		u:units = "meters s-1" ;
		u:grid = "fvcom_grid" ;
		u:type = "data" ;
	float v(time, siglay, nele) ;
		v:long_name = "Northward Water Velocity" ;
		v:units = "meters s-1" ;
		v:grid = "fvcom_grid" ;
		v:type = "data" ;
	float omega(time, siglev, node) ;
		omega:long_name = "Vertical Sigma Coordinate Velocity" ;
		omega:units = "s-1" ;
		omega:grid = "fvcom_grid" ;
		omega:type = "data" ;
	float ww(time, siglay, nele) ;
		ww:long_name = "Upward Water Velocity" ;
		ww:units = "meters s-1" ;
		ww:grid = "fvcom_grid" ;
		ww:type = "data" ;
	float ua(time, nele) ;
		ua:long_name = "Vertically Averaged x-velocity" ;
		ua:units = "meters s-1" ;
		ua:grid = "fvcom_grid" ;
		ua:type = "data" ;
	float va(time, nele) ;
		va:long_name = "Vertically Averaged y-velocity" ;
		va:units = "meters s-1" ;
		va:grid = "fvcom_grid" ;
		va:type = "data" ;
	float temp(time, siglay, node) ;
		temp:long_name = "temperature" ;
		temp:standard_name = "sea_water_temperature" ;
		temp:units = "degrees_C" ;
		temp:grid = "fvcom_grid" ;
		temp:coordinates = "x y" ;
		temp:type = "data" ;
	float salinity(time, siglay, node) ;
		salinity:long_name = "salinity" ;
		salinity:standard_name = "sea_water_salinity" ;
		salinity:units = "1e-3" ;
		salinity:grid = "fvcom_grid" ;
		salinity:coordinates = "x y" ;
		salinity:type = "data" ;

// global attributes:
		:title = "GDcoast case" ;
		:institution = "School for Marine Science and Technology" ;
		:source = "FVCOM_3.0" ;
		:Conventions = "CF-1.0" ;
		:CoordinateSystem = "Cartesian" ;
		:CoordinateProjection = "none: A recognized reference coordinate for projtion for PROJ4" ;
}
